library IEEE;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mipsFd is
	port (
        -- PORTAS ENTRADA
        CLK             : in STD_LOGIC;

        --UNIDADE DE CONTROLE
        MUX_PC_BEQ_JMP  : in STD_LOGIC;
        MUX_RT_RD       : in STD_LOGIC;
        HAB_ESCRITA_REG : in STD_LOGIC;

        HAB_LEITURA_MEM : in STD_LOGIC;
        HAB_ESCRITA_MEM : in STD_LOGIC;

        MUX_RT_IMM      : in STD_LOGIC;
        ULA_OP          : in STD_LOGIC_VECTOR(1 DOWNTO 0);
        MUX_ULA_MEM     : in STD_LOGIC;
        BEQ             : in STD_LOGIC;
        
        INST_OPCODE     : out STD_LOGIC_VECTOR(5 DOWNTO 0);   --OPCODE SAIDA
     


        --PLACA
        PC_RESET		: in STD_LOGIC;         


        -- DEBUG
        DEBUG_MEM_OUT			: out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_DADO_LIDO_1       : out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_DADO_LIDO_2       : out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_ULA_OUT			: out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_AUX_OP_OUT		: out STD_LOGIC_VECTOR(3 DOWNTO 0);
        DEBUG_AUX_HM            : out STD_LOGIC;
        DEBUG_ZERO_aux	        : out STD_LOGIC;
        DEBUG_MEM_W             : out STD_LOGIC_VECTOR(31 DOWNTO 0);
		  DEBUG_MEM_R				  : out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_DATA_MEM_ADDR     : out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_PC_OUT            : out STD_LOGIC_VECTOR(31 DOWNTO 0);
        DEBUG_PC4_BADD          : out STD_LOGIC_VECTOR(31 DOWNTO 0);
		  DEBUG_WRITE_REGISTER    : out STD_LOGIC_VECTOR(4 DOWNTO 0);
		  DEBUG_HAB_ESCRITA_REG	  : out STD_LOGIC;
		  DEBUG_WRITE_DATA    	  : out STD_LOGIC_VECTOR(31 DOWNTO 0);
		  DEBUG_SEL_ULA_MEM		  : out STD_LOGIC

    );

end entity;

architecture mipsFdArch of mipsFd is
    constant FOUR: STD_LOGIC_VECTOR(31 downto 0) := std_logic_vector(to_unsigned(4, 32));

    signal aux_pc_in            : STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
    signal aux_pc_out           : STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
    signal aux_mux_beq_out      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_mem_inst_out     : STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
    signal aux_som_pc_out       : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_banco_reg1_out   : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_banco_reg2_out   : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_extensor_out     : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_mux_rt_imm_out   : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_op               : STD_LOGIC_VECTOR(3 DOWNTO 0);
    signal aux_ula_out          : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_shifter32_out    : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_shifter26_out    : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_som_beq_out      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_ula_mem_out      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_ula_z            : STD_LOGIC;
    signal aux_mux_rt_rd_out    : STD_LOGIC_VECTOR(4 DOWNTO 0);
    signal aux_pc_reset         : STD_LOGIC := '0';

    signal aux_ifid_pc4         : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_ifid_inst        : STD_LOGIC_VECTOR(31 DOWNTO 0);
    
    
    signal aux_idex_wb          : STD_LOGIC_VECTOR(1 DOWNTO 0);
    signal aux_idex_m           : STD_LOGIC_VECTOR(2 DOWNTO 0);
    signal aux_idex_ex          : STD_LOGIC_VECTOR(3 DOWNTO 0);
    signal aux_idex_pc4         : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_idex_r1          : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_idex_r2          : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_idex_extend      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_idex_i16         : STD_LOGIC_VECTOR(4 DOWNTO 0);    
    signal aux_idex_i11         : STD_LOGIC_VECTOR(4 DOWNTO 0);
    

    signal aux_exmem_wb          : STD_LOGIC_VECTOR(1 DOWNTO 0);
    signal aux_exmem_m           : STD_LOGIC_VECTOR(2 DOWNTO 0);
    signal aux_exmem_som_beq     : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_exmem_z           : STD_LOGIC;
    signal aux_exmem_ular        : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_exmem_wd          : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_exmem_rtrd        : STD_LOGIC_VECTOR(4 DOWNTO 0);        

    signal aux_memwb_wb          : STD_LOGIC_VECTOR(1 DOWNTO 0);
    signal aux_memwb_data_mem_r  : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_memwb_end_mem     : STD_LOGIC_VECTOR(31 DOWNTO 0);
    signal aux_memwb_rtrd        : STD_LOGIC_VECTOR(4 DOWNTO 0);

    signal pc_src                : STD_LOGIC;
    signal aux_data_mem_r        : STD_LOGIC_VECTOR(31 DOWNTO 0);

--    signal terra                 : STD_LOGIC := '0';

begin
    IFID            : entity work.registradorGenerico 
                      generic map(larguraDados => 64) 
                      port map (
                            DIN(31 DOWNTO 0) =>  aux_mem_inst_out,
                            DIN(63 DOWNTO 32)  =>  aux_som_pc_out,
                            DOUT(31 DOWNTO 0) =>  aux_ifid_inst,  
                            DOUT(63 DOWNTO 32)=>  aux_ifid_pc4,
                            ENABLE => '1', 
                            CLK => CLK, 
                            RST => '0'
                      );


    IDEX            : entity work.registradorGenerico generic map(larguraDados => 147) port map(
        DIN(4 DOWNTO 0)     => aux_ifid_inst(15 DOWNTO 11),
        DIN(9 DOWNTO 5)     => aux_ifid_inst(20 DOWNTO 16),
        DIN(41 DOWNTO 10)   => aux_extensor_out,
        DIN(73 DOWNTO 42)   => aux_banco_reg2_out,
        DIN(105 DOWNTO 74)  => aux_banco_reg1_out, 
        DIN(137 DOWNTO 106) => aux_ifid_pc4,
        DIN(141 DOWNTO 138) => MUX_RT_RD & ULA_OP & MUX_RT_IMM,        
        DIN(144 DOWNTO 142) => BEQ & HAB_LEITURA_MEM & HAB_ESCRITA_MEM,
        DIN(146 DOWNTO 145) => HAB_ESCRITA_REG & MUX_ULA_MEM,

        DOUT(146 DOWNTO 145)=> aux_idex_wb,
        DOUT(144 DOWNTO 142)=> aux_idex_m,
        DOUT(141 DOWNTO 138)=> aux_idex_ex,
        DOUT(137 DOWNTO 106)=> aux_idex_pc4,
        DOUT(105 DOWNTO 74) => aux_idex_r1,
        DOUT(73 DOWNTO 42)  => aux_idex_r2,
        DOUT(41 DOWNTO 10)  => aux_idex_extend,
        DOUT(9 DOWNTO 5)    => aux_idex_i16,
        DOUT(4 DOWNTO 0)    => aux_idex_i11,

        ENABLE => '1',
        CLK => CLK,
        RST => '0'
    );

    EXMEM           : entity work.registradorGenerico generic map(larguraDados => 107) port map(
        DIN(4 DOWNTO 0)     => aux_mux_rt_rd_out,
        DIN(36 DOWNTO 5)    => aux_idex_r2,
        DIN(68 DOWNTO 37)   => aux_ula_out,
        DIN(69)             => aux_ula_z,
        DIN(101 DOWNTO 70)  => aux_som_beq_out,
        DIN(104 DOWNTO 102) => aux_idex_m,
        DIN(106 DOWNTO 105) => aux_idex_wb,

        DOUT(4 DOWNTO 0)    => aux_exmem_rtrd,
        DOUT(36 DOWNTO 5)   => aux_exmem_wd,
        DOUT(68 DOWNTO 37)  => aux_exmem_ular,
        DOUT(69)            => aux_exmem_z,
        DOUT(101 DOWNTO 70) => aux_exmem_som_beq,
        DOUT(104 DOWNTO 102)=> aux_exmem_m,
        DOUT(106 DOWNTO 105)=> aux_exmem_wb,
		  ENABLE => '1',
        CLK => CLK,
        RST => '0'
    );

    MEMWB            : entity work.registradorGenerico generic map(larguraDados => 71) port map (
        DIN(4 DOWNTO 0)     => aux_exmem_rtrd,
        DIN(36 DOWNTO 5)    => aux_exmem_ular,
        DIN(68 DOWNTO 37)   => aux_data_mem_r,
        DIN(70 DOWNTO 69)   => aux_exmem_wb,

        DOUT(4 DOWNTO 0)     => aux_memwb_rtrd,
        DOUT(36 DOWNTO 5)    => aux_memwb_end_mem,
        DOUT(68 DOWNTO 37)   => aux_memwb_data_mem_r,
        DOUT(70 DOWNTO 69)   => aux_memwb_wb,
		  ENABLE => '1',
        CLK => CLK,
        RST => '0'
    );

    memoriaDeDados  : entity work.memoriaAll port map (
        CLK => CLK, END_MEM => aux_exmem_ular, DATA_MEM_W => aux_exmem_wd, RD => aux_exmem_m(1), WR => aux_exmem_m(0), 
        DATA_MEM_R => aux_data_mem_r, HM => DEBUG_AUX_HM
    );

	PC				: entity work.registradorGenerico port map(DIN => aux_pc_in, DOUT => aux_pc_out, ENABLE => '1', CLK => CLK, RST => aux_pc_reset);
    memoriaDeInst   : entity work.memoriaDeInst port map(ADDR => to_integer(unsigned(aux_pc_out(31 DOWNTO 2))), CLK => CLK, Q => aux_mem_inst_out);
    bancoReg        : entity work.bancoRegistradores port map(
        HAB_ESCRITA_REG => aux_memwb_wb(1), CLK => CLK,
        END1 => aux_ifid_inst(25 DOWNTO 21), END2 => aux_ifid_inst(20 DOWNTO 16), END3 => aux_memwb_rtrd,
        DADO_W_REG3 => aux_ula_mem_out,
        DADO_R_REG1 => aux_banco_reg1_out, DADO_R_REG2 => aux_banco_reg2_out
    );

    ula             : entity work.ulaMips port map(
        A => aux_idex_r1, B => aux_mux_rt_imm_out, SEL => aux_op(1 DOWNTO 0), INVERTE_A => aux_op(3), INVERTE_B => aux_op(2), CIN => aux_op(2),
        R => aux_ula_out, ZERO => aux_ula_z
    ); 
	 
    ucUla           : entity work.ulaUc port map(FUNCT => aux_idex_extend(5 DOWNTO 0), ULA_OP => aux_idex_ex(2 DOWNTO 1), Q => aux_op);

    somadorPc       : entity work.somador port map(A => FOUR, B => aux_pc_out, Q => aux_som_pc_out);
    somadorBeq      : entity work.somador port map(A => aux_shifter32_out, B => aux_idex_pc4, Q => aux_som_beq_out);

    extensorSinal   : entity work.extensorSinal port map(A => aux_ifid_inst(15 DOWNTO 0), Q => aux_extensor_out); -- entra 16 sai 32

    shifter2_26     : entity work.shifterLeft2 port map(A => "000000" & aux_ifid_inst(25 DOWNTO 0), Q => aux_shifter26_out);
    shifter2_32     : entity work.shifterLeft2 port map(A => aux_idex_extend, Q => aux_shifter32_out);
    
    muxPc           : entity work.mux4 port map(A => aux_som_pc_out, B => aux_exmem_som_beq, C => aux_som_pc_out(31 DOWNTO 28) & aux_shifter26_out(27 DOWNTO 0), D => (others => '0'), SEL =>  MUX_PC_BEQ_JMP & pc_src, Q => aux_pc_in);

    muxRtRd         : entity work.mux2 generic map (data_len => 5) port map(A =>  aux_idex_i16, B =>  aux_idex_i11, SEL => aux_idex_ex(3), Q => aux_mux_rt_rd_out);
    muxRtImm        : entity work.mux2 port map(A => aux_idex_r2, B => aux_idex_extend, SEL => aux_idex_ex(0), Q => aux_mux_rt_imm_out);
    muxUlaMem       : entity work.mux2 port map(A => aux_memwb_data_mem_r, B => aux_memwb_end_mem, SEL => not aux_memwb_wb(0), Q => aux_ula_mem_out);     

    pc_src <= aux_exmem_m(2) and aux_exmem_z;
--    terra <= '0';

    --OPCODE SAIDA PRO FD
    INST_OPCODE <= aux_ifid_inst(31 downto 26);

    --ENTRADA DA PLACA
    aux_pc_reset <= PC_RESET;


    --DEBUG
    DEBUG_MEM_OUT			 <= aux_ifid_inst;
    DEBUG_DADO_LIDO_1        <= aux_idex_r1;
    DEBUG_DADO_LIDO_2        <= aux_idex_r2;
    DEBUG_ULA_OUT			 <= aux_exmem_ular;
    DEBUG_AUX_OP_OUT		 	<= aux_op;
--    DEBUG_AUX_HM             <= terra;--
    DEBUG_ZERO_aux	        <= aux_exmem_z;
    DEBUG_MEM_W              <= aux_exmem_wd;
    DEBUG_DATA_MEM_ADDR      <= aux_exmem_ular;
    DEBUG_PC_OUT             <= aux_pc_out;
    DEBUG_PC4_BADD           <= aux_exmem_som_beq;
	 DEBUG_MEM_R				  <= aux_memwb_data_mem_r;
	 DEBUG_WRITE_REGISTER	  <= aux_memwb_rtrd;
	 DEBUG_HAB_ESCRITA_REG    <= aux_memwb_wb(1);
	 DEBUG_WRITE_DATA			  <= aux_ula_mem_out;
	 DEBUG_SEL_ULA_MEM			<= aux_memwb_wb(0);
	 
end architecture;
